library ieee;
use ieee.std_logic_1164.all;

entity Cadeado5 is
	port(
		SW: in std_logic_vector(0 downto 0);
		Z: out std_logic
   );
end Cadeado5;

architecture behavior of Cadeado5 is
begin

end;
